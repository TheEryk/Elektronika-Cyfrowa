----------------------------------------------------------------------------------
-- Company: CCE
-- Engineer: Kropidlowski Marek
-- 
-- Create Date:    10:40:02 14/02/2015 
-- Description: generator przebiegow prostokatnych sterowany Bluetooth
--      wersja Nexys2
--      zakres: 0 .. 66 000 000 Hz
--      wypelnienie: 50%
--      rozdzielczosc regulacji: 1Hz
--      ustawienie warto�ci: liczba w Hz + znak 's'  (x"73")
--      
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity gen66_BT is
    Generic (pmodName : string := "JB");
    Port ( clk_50MHz : in  STD_LOGIC;
           -- led_test : out std_logic_vector(7 downto 0);
           -- sys_bus: bt_CTS,bt_RTS,bt_rst,bt_pair,bt_tx,bt_rx
           sys_bus : inout std_logic_vector(5 downto 0); -- LOC free
           f_out : out STD_LOGIC);
end gen66_BT;

----------------------------------------------------------------------------------
----------------------------------------------------------------------------------









----------------------------------------------------------------------------------
-- Module Name:    dds_gen - Behavioral 
-- Description: generator DDS, liczy wg wzoru:
--              fout = M * fclk/2^N
--   M - wspol. skalujacy akumulator fazy
--   N - szerokosc akumulatora fazy
--   sw - zadawana f, w Hz
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity dds_gen_v2 is
    Port ( clk : in  STD_LOGIC;
           sw : in  STD_LOGIC_VECTOR (25 downto 0);
           fout : out  STD_LOGIC);
end dds_gen_v2;

architecture Behavioral of dds_gen_v2 is
constant N: positive:=58; 
constant fclk: real:=200.0E6;
constant S: real:=(2.0**N)/fclk;
signal M, phase, phase_next: std_logic_vector(N-1 downto 0):=(others=>'0');

begin

M_calk: process(sw)
begin
  M <= sw * conv_std_logic_vector(integer(S),32);  
end process;

phase_acc: process(clk)
begin
  if rising_edge(clk) then
    phase_next <= phase;
  end if;
end process;

phase <= phase_next + M;
fout <= phase_next(N-1);

end Behavioral;

---------------------------------------------------------------------
--Device: xc3s500e-4fg320
--
-- Module dcm_4x
-- Generated by Xilinx Architecture Wizard
-- Written for synthesis tool: XST
-- Period Jitter (unit interval) for block DCM_SP_INST = 0.14 UI
-- Period Jitter (Peak-to-Peak) for block DCM_SP_INST = 0.70 ns
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;
library UNISIM;
use UNISIM.Vcomponents.ALL;

entity dcm_4x is
   port ( CLKIN_IN        : in    std_logic; 
          RST_IN          : in    std_logic; 
          CLKFX_OUT       : out   std_logic; 
          CLKIN_IBUFG_OUT : out   std_logic; 
          CLK0_OUT        : out   std_logic; 
          LOCKED_OUT      : out   std_logic);
end dcm_4x;

architecture BEHAVIORAL of dcm_4x is
   signal CLKFB_IN        : std_logic;
   signal CLKFX_BUF       : std_logic;
   signal CLKIN_IBUFG     : std_logic;
   signal CLK0_BUF        : std_logic;
   signal GND_BIT         : std_logic;
begin
   GND_BIT <= '0';
   CLKIN_IBUFG_OUT <= CLKIN_IBUFG;
   CLK0_OUT <= CLKFB_IN;
   CLKFX_BUFG_INST : BUFG
      port map (I=>CLKFX_BUF,
                O=>CLKFX_OUT);
   
--   CLKIN_IBUFG_INST : IBUFG
--      port map (I=>CLKIN_IN,
--                O=>CLKIN_IBUFG);
   
   CLK0_BUFG_INST : BUFG
      port map (I=>CLK0_BUF,
                O=>CLKFB_IN);
   
   DCM_SP_INST : DCM_SP
   generic map( CLK_FEEDBACK => "1X",
            CLKDV_DIVIDE => 2.0,
            CLKFX_DIVIDE => 1,
            CLKFX_MULTIPLY => 4,
            CLKIN_DIVIDE_BY_2 => FALSE,
            CLKIN_PERIOD => 20.000,
            CLKOUT_PHASE_SHIFT => "NONE",
            DESKEW_ADJUST => "SYSTEM_SYNCHRONOUS",
            DFS_FREQUENCY_MODE => "LOW",
            DLL_FREQUENCY_MODE => "LOW",
            DUTY_CYCLE_CORRECTION => TRUE,
            FACTORY_JF => x"C080",
            PHASE_SHIFT => 0,
            STARTUP_WAIT => FALSE)
      port map (CLKFB=>CLKFB_IN,
                CLKIN=>clkin_in, --CLKIN_IBUFG,
                DSSEN=>GND_BIT,
                PSCLK=>GND_BIT,
                PSEN=>GND_BIT,
                PSINCDEC=>GND_BIT,
                RST=>RST_IN,
                CLKDV=>open,
                CLKFX=>CLKFX_BUF,
                CLKFX180=>open,
                CLK0=>CLK0_BUF,
                CLK2X=>open,
                CLK2X180=>open,
                CLK90=>open,
                CLK180=>open,
                CLK270=>open,
                LOCKED=>LOCKED_OUT,
                PSDONE=>open,
                STATUS=>open);
   
end BEHAVIORAL;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
-- nexys2 bluetooth module
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library unisim;
use unisim.vcomponents.all;

entity Nx2_BT is
    Generic (pmodName : string := "JA");
    Port (
            -- system
            -- sys_bus: bt_CTS,bt_RTS,bt_rst,bt_pair,bt_tx,bt_rx
            sys_bus : inout std_logic_vector(5 downto 0); 
            -- user
            rx_bt : in std_logic; -- to BTM
            tx_bt : out std_logic -- from BTM
         );
end Nx2_BT;

architecture simple of Nx2_BT is
 ------------------------------------------------------------------------------
type pins_table is array(1 to 4) of string(1 to 23);
                                  -- jx4,jx3,jx8,jx7,jx9,jx10
constant pmod_table: pins_table := ("m15,l17,l16,k13,m14,m16", --A
                                    "t17,r15,r16,p17,t18,u18", --B
                                    "h16,g13,f14,h15,g16,j12", --C
                                    "p18,n18,k15,k14,j15,j14");--D
function address(x: string) return natural is
begin
    if x="JB" then return 2;
    elsif x="JC" then return 3;
    elsif x="JD" then return 4;
    else return 1;
    end if;
end function;

signal cts_i, rts_i, rst_i, pair_i, tx_i, rx_i: std_logic;

attribute keep: string;
attribute keep of sys_bus: signal is "TRUE";
attribute loc: string;
attribute loc of sys_bus: signal is pmod_table(address(pmodName));

begin
  -- bypass
rx_i <= rx_bt;
tx_bt <= tx_i;

  -- test
rst_i <= '0';
pair_i <= '0';
cts_i <= rts_i;

  -- fpga pins
obufcts: OBUF port map(I => cts_i, O => sys_bus(5));
ibufrts: IBUF port map(O => rts_i, I => sys_bus(4));
obufrst: OBUF port map(I => rst_i, O => sys_bus(3));
obufpair: OBUF port map(I => pair_i, O => sys_bus(2));
obufrx: OBUF port map(I => rx_i, O => sys_bus(0));
ibuftx: IBUF port map(O => tx_i, I => sys_bus(1));

end simple;
----------------------------------------------------------------------
-- BCD to binary conwerter
-- by HusTakocem 2014
--
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity bcd2bin is
  generic (N_digit: natural:=4);   -- bcd digit #
  port (Clock : in std_logic;
        Init : in std_logic;       -- initialise the BCD conversion
        BCD_in : in std_logic_vector((N_digit*4)-1 downto 0); -- BCD input
        Done : out std_logic;
        BIN_out : out std_logic_vector((N_digit*4)-1 downto 0) -- binary output
       );
end;

architecture behav of bcd2bin is
signal shift_reg: std_logic_vector(BCD_in'range):=(others=>'0');
signal reg_temp: std_logic_vector(BCD_in'range):=(others=>'0');
signal out_reg: std_logic_vector(BCD_in'range):=(others=>'0');
signal shift_cntr: std_logic_vector(7 downto 0):=(others=>'0');
signal ok: std_logic := '0';

function conversion(bcd: std_logic_vector(3 downto 0)) return std_logic_vector is
  variable slv: std_logic_vector(bcd'range);
  begin
    case bcd is
        when "0000" => slv := "0000";
        when "0001" => slv := "0001";
        when "0010" => slv := "0010";
        when "0011" => slv := "0011";
        when "0100" => slv := "0100";
        when "0101" => slv := "0101";
        when "0110" => slv := "0110";
        when "0111" => slv := "0111";
        when "1000" => slv := "0101";
        when "1001" => slv := "0110";
        when "1010" => slv := "0111";
        when "1011" => slv := "1000";
        when "1100" => slv := "1001";
        when "1101" => slv := "1010";
        when "1110" => slv := "1011";
        when "1111" => slv := "1100";
        when others => slv := (others => '-');
    end case;
    return slv;
  end function;
begin

reg_shitf: process(clock)
  begin
    if rising_edge(clock) then  
        if Init='1' then
            shift_reg <= '0' & BCD_in((N_digit*4)-1 downto 1);
            out_reg <= BCD_in(0) & conv_std_logic_vector(0,(N_digit*4)-1);
            shift_cntr <= (others => '0');
        elsif ok='0' then
            shift_reg <= '0' & reg_temp((N_digit*4)-1 downto 1);
            out_reg <= reg_temp(0) & out_reg((N_digit*4)-1 downto 1);
            shift_cntr <= shift_cntr + 1;
        else 
            shift_reg <= shift_reg;
            out_reg <= out_reg;
            shift_cntr <= shift_cntr;
        end if;
    end if;
end process;

reg_conversion: process(shift_reg)
begin
  for i in 1 to N_digit loop
    reg_temp((i*4)-1 downto (i*4)-4) <= conversion(shift_reg((i*4)-1 downto (i*4)-4));
  end loop;
end process;

ok <= '1' when shift_cntr=(N_digit*4)-1 else '0';
Done <= ok;
BIN_out <= out_reg;

end architecture;
-----------------------------------------------------------------------------------
-----------------------------------------------------------------------------------
-- Constant (K) Compact UART Receiver
--
-- Version : 1.10 
-- Version Date : 3rd December 2003
-- Reason : '--translate' directives changed to '--synthesis translate' directives
--
-- Version : 1.00
-- Version Date : 16th October 2002
--
-- Start of design entry : 16th October 2002
--
-- Ken Chapman
-- Xilinx Ltd
-- Benchmark House
-- 203 Brooklands Road
-- Weybridge
-- Surrey KT13 ORH
-- United Kingdom
--
-- chapman@xilinx.com
--
------------------------------------------------------------------------------------
--
-- NOTICE:
--
-- Copyright Xilinx, Inc. 2002.   This code may be contain portions patented by other 
-- third parties.  By providing this core as one possible implementation of a standard,
-- Xilinx is making no representation that the provided implementation of this standard 
-- is free from any claims of infringement by any third party.  Xilinx expressly 
-- disclaims any warranty with respect to the adequacy of the implementation, including 
-- but not limited to any warranty or representation that the implementation is free 
-- from claims of any third party.  Futhermore, Xilinx is providing this core as a 
-- courtesy to you and suggests that you contact all third parties to obtain the 
-- necessary rights to use this implementation.
--
------------------------------------------------------------------------------------
---
-- uart_rx
-- 
-- uart receiver with baudrate counter (main clock = 50MHz, terminal settings: 19200 8-N-1)
---
------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity uart_rx is
    Generic (BaudRate: positive := 19200);
    Port (        clk : in std_logic; -- 50MHz (Nexys2 - B8)
                   rx : in std_logic; -- serial_in (Nexys2 - U6)
             data_out : out std_logic_vector(7 downto 0); -- received char
          data_strobe : out std_logic); -- valid data
    end uart_rx;
------------------------------------------------------------------------------------
------------------------------------------------------------------------------------
--
-- Library declarations
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library unisim;
use unisim.vcomponents.all;
--
------------------------------------------------------------------------------------
--
-- Main Entity for KCUART_RX
--
entity kcuart_rx is
    Port (      serial_in : in std_logic;  
                 data_out : out std_logic_vector(7 downto 0);
              data_strobe : out std_logic;
             en_16_x_baud : in std_logic;
                      clk : in std_logic);
    end kcuart_rx;
--
------------------------------------------------------------------------------------
--
-- Start of Main Architecture for KCUART_RX
--	 
architecture low_level_definition of kcuart_rx is
--
------------------------------------------------------------------------------------
--
------------------------------------------------------------------------------------
--
-- Signals used in KCUART_RX
--
------------------------------------------------------------------------------------
--
signal sync_serial        : std_logic;
signal stop_bit           : std_logic;
signal data_int           : std_logic_vector(7 downto 0);
signal data_delay         : std_logic_vector(7 downto 0);
signal start_delay        : std_logic;
signal start_bit          : std_logic;
signal edge_delay         : std_logic;
signal start_edge         : std_logic;
signal decode_valid_char  : std_logic;
signal valid_char         : std_logic;
signal decode_purge       : std_logic;
signal purge              : std_logic;
signal valid_srl_delay    : std_logic_vector(8 downto 0);
signal valid_reg_delay    : std_logic_vector(8 downto 0);
signal decode_data_strobe : std_logic;
--
--
------------------------------------------------------------------------------------
--
-- Attributes to define LUT contents during implementation 
-- The information is repeated in the generic map for functional simulation--
--
------------------------------------------------------------------------------------
--
attribute INIT : string; 
attribute INIT of start_srl     : label is "0000";
attribute INIT of edge_srl      : label is "0000";
attribute INIT of valid_lut     : label is "0040";
attribute INIT of purge_lut     : label is "54";
attribute INIT of strobe_lut    : label is "8";
--
------------------------------------------------------------------------------------
--
-- Start of KCUART_RX circuit description
--
------------------------------------------------------------------------------------
--	
begin

  -- Synchronise input serial data to system clock

  sync_reg: FD
  port map ( D => serial_in,
             Q => sync_serial,
             C => clk);

  stop_reg: FD
  port map ( D => sync_serial,
             Q => stop_bit,
             C => clk);


  -- Data delays to capture data at 16 time baud rate
  -- Each SRL16E is followed by a flip-flop for best timing

  data_loop: for i in 0 to 7 generate
  begin

     lsbs: if i<7 generate
     --
     attribute INIT : string; 
     attribute INIT of delay15_srl : label is "0000"; 
     --
     begin

       delay15_srl: SRL16E
       --synthesis translate_off
       generic map (INIT => X"0000")
       --synthesis translate_on
       port map(   D => data_int(i+1),
                  CE => en_16_x_baud,
                 CLK => clk,
                  A0 => '0',
                  A1 => '1',
                  A2 => '1',
                  A3 => '1',
                   Q => data_delay(i) );

     end generate lsbs;

     msb: if i=7 generate
     --
     attribute INIT : string; 
     attribute INIT of delay15_srl : label is "0000"; 
     --
     begin

       delay15_srl: SRL16E
       --synthesis translate_off
       generic map (INIT => X"0000")
       --synthesis translate_on
       port map(   D => stop_bit,
                  CE => en_16_x_baud,
                 CLK => clk,
                  A0 => '0',
                  A1 => '1',
                  A2 => '1',
                  A3 => '1',
                   Q => data_delay(i) );

     end generate msb;

     data_reg: FDE
     port map ( D => data_delay(i),
                Q => data_int(i),
               CE => en_16_x_baud,
                C => clk);

  end generate data_loop;

  -- Assign internal signals to outputs

  data_out <= data_int;
 
  -- Data delays to capture start bit at 16 time baud rate

  start_srl: SRL16E
  --synthesis translate_off
  generic map (INIT => X"0000")
  --synthesis translate_on
  port map(   D => data_int(0),
             CE => en_16_x_baud,
            CLK => clk,
             A0 => '0',
             A1 => '1',
             A2 => '1',
             A3 => '1',
              Q => start_delay );

  start_reg: FDE
  port map ( D => start_delay,
             Q => start_bit,
            CE => en_16_x_baud,
             C => clk);


  -- Data delays to capture start bit leading edge at 16 time baud rate
  -- Delay ensures data is captured at mid-bit position

  edge_srl: SRL16E
  --synthesis translate_off
  generic map (INIT => X"0000")
  --synthesis translate_on
  port map(   D => start_bit,
             CE => en_16_x_baud,
            CLK => clk,
             A0 => '1',
             A1 => '0',
             A2 => '1',
             A3 => '0',
              Q => edge_delay );

  edge_reg: FDE
  port map ( D => edge_delay,
             Q => start_edge,
            CE => en_16_x_baud,
             C => clk);

  -- Detect a valid character 

  valid_lut: LUT4
  --synthesis translate_off
  generic map (INIT => X"0040")
  --synthesis translate_on
  port map( I0 => purge,
            I1 => stop_bit,
            I2 => start_edge,
            I3 => edge_delay,
             O => decode_valid_char );  

  valid_reg: FDE
  port map ( D => decode_valid_char,
             Q => valid_char,
            CE => en_16_x_baud,
             C => clk);

  -- Purge of data status 

  purge_lut: LUT3
  --synthesis translate_off
  generic map (INIT => X"54")
  --synthesis translate_on
  port map( I0 => valid_reg_delay(8),
            I1 => valid_char,
            I2 => purge,
             O => decode_purge );  

  purge_reg: FDE
  port map ( D => decode_purge,
             Q => purge,
            CE => en_16_x_baud,
             C => clk);

  -- Delay of valid_char pulse of length equivalent to the time taken 
  -- to purge data shift register of all data which has been used.
  -- Requires 9x16 + 8 delays which is achieved by packing of SRL16E with 
  -- up to 16 delays and utilising the dedicated flip flop in each stage.

  valid_loop: for i in 0 to 8 generate
  begin

     lsb: if i=0 generate
     --
     attribute INIT : string; 
     attribute INIT of delay15_srl : label is "0000"; 
     --
     begin

       delay15_srl: SRL16E
       --synthesis translate_off
       generic map (INIT => X"0000")
       --synthesis translate_on
       port map(   D => valid_char,
                  CE => en_16_x_baud,
                 CLK => clk,
                  A0 => '0',
                  A1 => '1',
                  A2 => '1',
                  A3 => '1',
                   Q => valid_srl_delay(i) );

     end generate lsb;

     msbs: if i>0 generate
     --
     attribute INIT : string; 
     attribute INIT of delay16_srl : label is "0000"; 
     --
     begin

       delay16_srl: SRL16E
       --synthesis translate_off
       generic map (INIT => X"0000")
       --synthesis translate_on
       port map(   D => valid_reg_delay(i-1),
                  CE => en_16_x_baud,
                 CLK => clk,
                  A0 => '1',
                  A1 => '1',
                  A2 => '1',
                  A3 => '1',
                   Q => valid_srl_delay(i) );

     end generate msbs;

     data_reg: FDE
     port map ( D => valid_srl_delay(i),
                Q => valid_reg_delay(i),
               CE => en_16_x_baud,
                C => clk);

  end generate valid_loop;

  -- Form data strobe

  strobe_lut: LUT2
  --synthesis translate_off
  generic map (INIT => X"8")
  --synthesis translate_on
  port map( I0 => valid_char,
            I1 => en_16_x_baud,
             O => decode_data_strobe );

  strobe_reg: FD
  port map ( D => decode_data_strobe,
             Q => data_strobe,
             C => clk);

end low_level_definition;

--------------------------------------------------------------------

architecture mixed of uart_rx is
-- baud_count = fclk/(baud_rate * 16)
constant baud_val: natural := 50E6/BaudRate/16;

    component kcuart_rx is
    Port (    serial_in : in std_logic;  
               data_out : out std_logic_vector(7 downto 0);
            data_strobe : out std_logic;
           en_16_x_baud : in std_logic;
                    clk : in std_logic);
    end component;

    -- UART signals
    signal baud_count   : std_logic_vector (8 downto 0):=(others=>'0');
    signal en_16_x_baud : std_logic:='0';

begin
    
    baudgen: process (clk)
    begin  
    if (clk'event and clk = '1') then
        if (baud_count = baud_val)then
                baud_count <= (others=>'0');
                en_16_x_baud <= '1';
        else
                baud_count <= baud_count + 1;
                en_16_x_baud <= '0';
        end if;
    end if;
    end process;

    receiver: kcuart_rx
    port map (rx, data_out, data_strobe, en_16_x_baud, clk);

end architecture;
-------------------------------------------------------------------------------------
-- gen_ctrl
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity gen_ctrl is
  port (clk : in std_logic;
        strobe : in std_logic;
        data : in std_logic_vector(7 downto 0);
        init : out std_logic;
        bcd : out std_logic_vector(31 downto 0)); -- 8 digit
end entity;

architecture fsm of gen_ctrl is
constant Set: std_logic_vector(7 downto 0):=x"73"; -- char s
type digit_array is array (8 downto 0) of std_logic_vector(3 downto 0); -- 8 digit + command
type fsm_state is (idle,reg_reset,get_char,set_out);
signal state,xstate: fsm_state;
signal bcd_reg : digit_array := (others=>x"0");
signal init_string : boolean;
signal init_i, reset : std_logic;

begin

fsm: process(state,strobe,init_string)
begin
    case state is
        when idle => if strobe='1' then xstate <= get_char; else xstate <= idle; end if;
        when get_char => if init_string then xstate <= set_out; else xstate <= idle; end if;
        when set_out => xstate <= reg_reset;
        when reg_reset => xstate <= idle;
        when others => xstate <= idle;
    end case;
end process; 

fsm_reg: process(clk)
begin
    if rising_edge(clk) then
        state <= xstate;
    end if;
end process;

get_data:process(clk)
begin
    if rising_edge(clk) then
      if reset='1' then
        bcd_reg <= (others=>x"0");
      elsif strobe='1' then
        bcd_reg <= bcd_reg(7 downto 0) & data(3 downto 0);
      end if;
    end if;
end process;

init_string <= true when data=Set else false;
init_i <= '1' when state = set_out else '0';
reset <= '1' when state = reg_reset else '0';
init <= init_i;
bcd <= bcd_reg(8) & bcd_reg(7) & bcd_reg(6) & bcd_reg(5) & bcd_reg(4) & bcd_reg(3) & bcd_reg(2) & bcd_reg(1);

end architecture;
-------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------
architecture mix of gen66_BT is

constant N_gen: natural := 26;
signal bcd : std_logic_vector(31 downto 0);
signal bin_freq : std_logic_vector(31 downto 0);
signal clk_4x, clk_slow_en, btn_up_en, btn_shift_en, btn_down_en: std_logic;
signal serial_data, bypass, valid_data, init, done : std_logic;
signal clk_50MHz_dcm: std_logic;
signal data_from_BT : std_logic_vector(7 downto 0);

begin

dds: entity work.dds_gen_v2
    port map(clk_4x,bin_freq(N_gen-1 downto 0),f_out);
    
mul4: entity work.dcm_4x
    port map(CLKIN_IN=>clk_50MHz,RST_IN=>'0',CLKFX_OUT=>clk_4x, CLK0_OUT=>clk_50MHz_dcm);
    
BT: entity work.Nx2_BT
    generic map(pmodName => pmodName)
    Port map(sys_bus => sys_bus,rx_bt => bypass,tx_bt => serial_data);
    bypass <= serial_data; -- echo

uart: entity work.uart_rx
    Generic map (BaudRate => 19200)
    Port map( clk => clk_50MHz_dcm, rx => serial_data, 
              data_out => data_from_bt, data_strobe => valid_data);
    
bcd_conv: entity work.bcd2bin
    generic map (N_digit => 8)   -- bcd digit #
    port map (Clock => clk_50MHz_dcm,Init => init,BCD_in => bcd,Done => done,BIN_out => bin_freq);
        
ctrl: entity work.gen_ctrl
    port map (clk => clk_50MHz_dcm,strobe => valid_data,data => data_from_bt,init => init,
              bcd => bcd); -- out std_logic_vector(31 downto 0)); -- 8 digit

end architecture;